`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/15/2024 07:44:43 PM
// Design Name: 
// Module Name: reg_file
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module reg_file(
    input wire CLK,
    input wire RegWrite1,        // Write enable for the first register
    input wire RegWrite2,        // Write enable for the second register
    input wire [2:0] srcA,       // Source register A address
    input wire [2:0] srcB,       // Source register B address
    input wire [2:0] writeReg1,  // First destination register address
    input wire [2:0] writeReg2,  // Second destination register address
    input wire [9:0] writeValue1,// Value to write to the first register
    input wire [9:0] writeValue2,// Value to write to the second register
    output [9:0] ReadA,          // Data read from source A
    output [9:0] ReadB           // Data read from source B
);

    wire [7:0] writeEnable1, writeEnable2;  // One-hot write enable signals
    wire [9:0] registers [7:0];             // 8 registers, each 10 bits wide

    // One-hot Write Enable signals generated by decoders
    decoder_3to8 decoder1 (
        .addr(writeReg1),
        .enable(RegWrite1),
        .out(writeEnable1)
    );

    decoder_3to8 decoder2 (
        .addr(writeReg2),
        .enable(RegWrite2),
        .out(writeEnable2)
    );

    // Instantiate 8 DFF modules for each register
    genvar i;
    generate
        for (i = 0; i < 8; i = i + 1) begin : reg_loop
            dff_10bit dff (
                .CLK(CLK),
                .D(writeEnable1[i] ? writeValue1 : writeValue2), // Write Value Priority
                .enable(writeEnable1[i] | writeEnable2[i]),      // Enable condition
                .Q(registers[i])
            );
        end
    endgenerate

    // Read outputs using multiplexers
    mux8x1 muxA (
        .reg0(registers[0]), .reg1(registers[1]), .reg2(registers[2]),
        .reg3(registers[3]), .reg4(registers[4]), .reg5(registers[5]),
        .reg6(registers[6]), .reg7(registers[7]),
        .sel(srcA),
        .out(ReadA)
    );

    mux8x1 muxB (
        .reg0(registers[0]), .reg1(registers[1]), .reg2(registers[2]),
        .reg3(registers[3]), .reg4(registers[4]), .reg5(registers[5]),
        .reg6(registers[6]), .reg7(registers[7]),
        .sel(srcB),
        .out(ReadB)
    );

endmodule
